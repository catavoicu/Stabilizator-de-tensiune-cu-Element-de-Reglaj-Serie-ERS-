** Profile: "SCHEMATIC1-Sarcina"  [ C:\Users\catav\OneDrive - Universitatea Politehnica Bucuresti\Desktop\P1\p1_voicu_catalin-pspicefiles\schematic1\sarcina.sim ] 

** Creating circuit file "Sarcina.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "c:/cadence/orcadx_24.1/tools/capture/library/p1/bc846b.lib" 
.LIB "c:/cadence/orcadx_24.1/tools/capture/library/p1/bc856b.lib" 
.LIB "c:/cadence/orcadx_24.1/tools/capture/library/p1/bzx84c10.lib" 
.LIB "c:/cadence/orcadx_24.1/tools/capture/library/p1/mjd31cg.lib" 
* From [PSPICE NETLIST] section of C:\Users\catav\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM Rload 10 100 0.1 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
